`timescale 1ns / 1ps

module Main(
    input Clk,
    input [7:0] N,
    input Start,
    output Salida,
	 output [7:0] Displays, Segmentos
    );
    
    wire a1_,a2_,a3_,a4_,a5_,a6_,a7_;
    wire [7:0] A_,E_,K_,Sal;
	 wire P;
    
    Data_path U1 (
    .clk(Clk),
    .n(N),
    .a1(a1_),
    .a2(a2_),
    .a3(a3_),
    .a4(a4_),
    .a5(a5_),
    .a6(a6_),
    .a7(a7_),
    .A(A_),
    .P(Salida),
	 .Sal(Sal),
    .K(K_),
    .E(E_)
    
    );
    FSM U2 (
    
    .clk(Clk),
    .start(Start),
    .A(A_),
    .E(E_),
    .K(K_),
    .a1(a1_),
    .a2(a2_),
    .a3(a3_),
    .a4(a4_),
    .a5(a5_),
    .a6(a6_),
    .a7(a7_) 
    );
	 
	 Multiplexor U3(
    .Clk(Clk), 
    .Displays(Displays), 
    .Segmentos(Segmentos), 
    .Sal(Sal), 
	 .Salida(Salida)
    );
	 

endmodule